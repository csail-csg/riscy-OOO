import Types::*;

Addr bootRomBaseAddr = 64'h00001000;
Addr msipBaseAddr    = 64'h02000000;
Addr mtimcmpBaseAddr = 64'h02004000;
Addr mtimeBaseAddr   = 64'h0200bff8;
Addr mainMemBaseAddr = 64'h80000000;

