
// Copyright (c) 2017 Massachusetts Institute of Technology
// 
// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:
// 
// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.
// 
// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import Types::*;
import ProcTypes::*;
import Core::*;
import CrossBar::*;
import Vector::*;
import GetPut::*;

module mkIPIConnect#(Vector#(CoreNum, CoreIPI) ipi)(Empty);
    Vector#(CoreNum, Get#(CoreId)) src = ?;
    Vector#(CoreNum, Put#(void)) dst = ?;
    for(Integer i = 0; i < valueof(CoreNum); i = i+1) begin
        src[i] = toGet(ipi[i].sendIPI);
        dst[i] = (interface Put;
            method Action put(void x);
                ipi[i].recvIPI;
            endmethod
        endinterface);
    end

    function XBarDstInfo#(CoreId, void) getDst(CoreId srcIdx, CoreId srcData);
        return XBarDstInfo {idx: srcData, data: ?};
    endfunction
    mkXBar(getDst, src, dst);
endmodule
